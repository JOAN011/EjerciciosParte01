----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:59:17 07/11/2022 
-- Design Name: 
-- Module Name:    Registro_Paralelo - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Registro_Paralelo is
    Port ( D : in  STD_LOGIC_VECTOR (0 to 7);
           clk : in  STD_LOGIC;
           Q : out  STD_LOGIC_VECTOR (0 to 7));
end Registro_Paralelo;

architecture Behavioral of Registro_Paralelo is
begin
	process (clk) begin
	if (clk' event and clk = '1') then
		Q	<= D;
	end if;
	end process;
end Behavioral;

